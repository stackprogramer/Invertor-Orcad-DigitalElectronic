** Profile: "SCHEMATIC1-t"  [ F:\Users\ROOT\Documents\orcad\elecdigital\problem1\p1-schematic1-t.sim ] 

** Creating circuit file "p1-schematic1-t.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of F:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1s 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\p1-SCHEMATIC1.net" 


.END
