** Profile: "SCHEMATIC1-t"  [ F:\Users\ROOT\Documents\orcad\elecdigital\problem1 - asli\p2-schematic1-t.sim ] 

** Creating circuit file "p2-schematic1-t.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\p2.lib" 
* From [PSPICE NETLIST] section of F:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 .01 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\p2-SCHEMATIC1.net" 


.END
